module top_module(
    output zero
);
    assign zero=0;
endmodule

