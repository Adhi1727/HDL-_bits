module top_module(
    input clk,
    input areset,    
    input in,
    output out);

    parameter A=0;
    parameter B=1; 
    reg state, next_state;

    always @(*) begin
        case(state)
            A:if(in==0)
                next_state=B;
            else 
                next_state=A;
            B:if(in==0)
                next_state=A;
            else
                next_state=B;
        endcase
    end

    always @(posedge clk, posedge areset) begin
        if(areset)
            state<=B;
        else
            state<=next_state;
    end
            
    assign out = (state==B);
                
endmodule

